module tb();

    initial begin
        $hello;
    end

endmodule
